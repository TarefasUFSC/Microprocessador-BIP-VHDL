ROM_INTEL_SREG_inst : ROM_INTEL_SREG PORT MAP (
		address	 => address_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
